`timescale 1 ns / 100 ps

/*
	register file implemented based on the description 
	provided in Computer Organization and Design, 5th
*/

module register_file()


endmodule
